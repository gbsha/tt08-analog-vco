** sch_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_stage_half.sch
.subckt vco_stage_half VDD VSS Vin Vb Vd Vout Vs Vbuf
*.PININFO VDD:B VSS:B Vin:I Vb:I Vd:I Vout:O Vs:O Vbuf:O
XM7 Vout Vd VDD VDD sky130_fd_pr__pfet_01v8 L=2 W=4 nf=2 m=1
XM3 Vout Vb VDD VDD sky130_fd_pr__pfet_01v8 L=2 W=4 nf=2 m=1
XM1 Vout Vin Vs VSS sky130_fd_pr__nfet_01v8 L=2 W=4 nf=2 m=1
x1 VDD VSS Vout Vbuf vco_buffer
XM8 VSS Vout VSS VSS sky130_fd_pr__nfet_01v8 L=11 W=11 nf=1 m=1
.ends

* expanding   symbol:  vco_buffer.sym # of pins=4
** sym_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_buffer.sym
** sch_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_buffer.sch
.subckt vco_buffer VDD VSS Vin Vout
*.PININFO VDD:B VSS:B Vin:I Vout:O
x1 VDD Vin net1 VSS vco_inverter
x2 VDD net1 Vout VSS vco_inverter
.ends


* expanding   symbol:  vco_inverter.sym # of pins=4
** sym_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_inverter.sym
** sch_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_inverter.sch
.subckt vco_inverter VDD Vin Vout VSS
*.PININFO VDD:B VSS:B Vin:I Vout:O
XM1 Vout Vin VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
