magic
tech sky130A
magscale 1 2
timestamp 1725469944
<< locali >>
rect 1430 3200 4720 3250
rect 1430 3090 1690 3200
rect 4660 3090 4720 3200
rect 1430 2860 4720 3090
rect 1430 2240 2060 2860
rect 3480 2240 4720 2860
rect 1430 1330 1850 2240
rect 3650 1330 4720 2240
rect 1430 1140 4720 1330
rect 1430 400 2080 1140
rect 3650 1130 4720 1140
rect 4480 400 4720 1130
rect 1430 -2310 1990 240
rect 4500 -2310 4720 230
rect 1430 -2580 4720 -2310
rect 1430 -2620 2710 -2580
rect 3820 -2620 4720 -2580
rect 1430 -3360 2680 -2620
rect 3850 -3360 4720 -2620
rect 1430 -3390 4720 -3360
rect 1430 -3840 4730 -3390
rect 1430 -3970 1780 -3840
rect 4370 -3970 4730 -3840
rect 1430 -4000 4730 -3970
<< viali >>
rect 1690 3090 4660 3200
rect 1780 -3970 4370 -3840
<< metal1 >>
rect 1430 3200 4720 3250
rect 1430 3090 1690 3200
rect 4660 3090 4720 3200
rect 1430 3050 4720 3090
rect 2010 2700 2020 2900
rect 2230 2700 2240 2900
rect 2010 2090 2020 2290
rect 2220 2090 2230 2290
rect 3300 2090 4330 2290
rect 2010 1500 2020 1700
rect 2220 1500 2230 1700
rect 1430 1440 1630 1500
rect 1430 1370 4590 1440
rect 1430 1300 1630 1370
rect 1430 210 1690 410
rect 1890 350 1900 410
rect 2110 350 2170 980
rect 2370 490 2470 1370
rect 2600 580 2610 980
rect 2680 580 2690 980
rect 2840 500 2940 1370
rect 3470 1210 4720 1290
rect 3120 350 3180 980
rect 3360 350 3420 980
rect 3640 500 3750 1210
rect 3850 580 3860 980
rect 3930 580 3940 980
rect 4090 500 4200 1210
rect 4520 1090 4720 1210
rect 4370 350 4430 980
rect 1890 270 4640 350
rect 1890 210 1900 270
rect 2070 -2080 2080 20
rect 2150 -2080 2160 20
rect 3080 -2220 3310 270
rect 4340 -2090 4350 20
rect 4410 -2090 4420 20
rect 1430 -2400 1630 -2360
rect 1430 -2520 4720 -2400
rect 1430 -2560 1630 -2520
rect 2730 -3500 2790 -2720
rect 3000 -3190 3090 -2520
rect 3220 -3120 3230 -2720
rect 3300 -3120 3310 -2720
rect 3450 -3200 3540 -2520
rect 3740 -3500 3800 -2720
rect 4520 -3500 4720 -3430
rect 2730 -3560 4720 -3500
rect 4520 -3630 4720 -3560
rect 1430 -3840 4730 -3800
rect 1430 -3970 1780 -3840
rect 4370 -3970 4730 -3840
rect 1430 -4000 4730 -3970
<< via1 >>
rect 1690 3090 4660 3200
rect 2020 2700 2230 2900
rect 2020 2090 2220 2290
rect 2020 1500 2220 1700
rect 1690 210 1890 410
rect 2610 580 2680 980
rect 3860 580 3930 980
rect 2080 -2080 2150 20
rect 4350 -2090 4410 20
rect 3230 -3120 3300 -2720
rect 1780 -3970 4370 -3840
<< metal2 >>
rect 1630 3210 3950 3250
rect 1630 3200 4660 3210
rect 1630 3090 1690 3200
rect 1630 3080 4660 3090
rect 1630 3050 3950 3080
rect 2020 2900 2230 3050
rect 2020 2690 2230 2700
rect 2020 2290 2220 2300
rect 2020 2080 2220 2090
rect 2020 1700 2220 1710
rect 2020 1490 2220 1500
rect 1690 410 1890 420
rect 1690 200 1890 210
rect 2090 30 2150 1490
rect 2620 990 2670 3050
rect 3870 990 3920 3050
rect 2610 980 2680 990
rect 2610 570 2680 580
rect 3860 980 3930 990
rect 3860 570 3930 580
rect 2080 20 2150 30
rect 2080 -2090 2150 -2080
rect 2090 -3800 2150 -2090
rect 4350 20 4410 60
rect 3230 -2720 3300 -2710
rect 3230 -3130 3300 -3120
rect 4350 -3800 4410 -2090
rect 1750 -3840 4430 -3800
rect 1750 -3970 1780 -3840
rect 4370 -3970 4430 -3840
rect 1750 -4000 4430 -3970
<< via2 >>
rect 2020 2090 2220 2290
rect 1690 210 1890 410
rect 3230 -3120 3300 -2720
<< metal3 >>
rect 2010 2290 2230 2295
rect 1710 2090 2020 2290
rect 2220 2090 2230 2290
rect 1710 415 1850 2090
rect 2010 2085 2230 2090
rect 1680 410 1900 415
rect 1680 210 1690 410
rect 1890 210 1900 410
rect 1680 205 1900 210
rect 1710 -2870 1850 205
rect 3220 -2720 3310 -2715
rect 3220 -2870 3230 -2720
rect 1710 -2970 3230 -2870
rect 3220 -3120 3230 -2970
rect 3300 -3120 3310 -2720
rect 3220 -3125 3310 -3120
use vco_buffer  vco_buffer_0
timestamp 1725445236
transform 1 0 2020 0 1 1510
box 0 -10 1480 1390
use sky130_fd_pr__nfet_01v8_XVWV9B  XM1
timestamp 1725469944
transform 1 0 3265 0 1 -2920
box -625 -410 625 410
use sky130_fd_pr__pfet_01v8_GJP7VV  XM3
timestamp 1725457726
transform 1 0 2645 0 1 779
box -625 -419 625 419
use sky130_fd_pr__pfet_01v8_GJP7VV  XM7
timestamp 1725457726
transform 1 0 3895 0 1 779
box -625 -419 625 419
use sky130_fd_pr__nfet_01v8_APRB2X  XM8
timestamp 1725457726
transform 1 0 3246 0 1 -1040
box -1296 -1310 1296 1310
<< labels >>
flabel metal1 1430 3050 1630 3250 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1430 1300 1630 1500 0 FreeSans 256 0 0 0 Vb
port 3 nsew
flabel metal1 1430 210 1630 410 0 FreeSans 256 0 0 0 Vout
port 5 nsew
flabel metal1 4520 1090 4720 1290 0 FreeSans 256 0 0 0 Vd
port 4 nsew
flabel metal1 4130 2090 4330 2290 0 FreeSans 256 0 0 0 Vbuf
port 7 nsew
flabel metal1 1430 -2560 1630 -2360 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 4520 -3630 4720 -3430 0 FreeSans 256 0 0 0 Vs
port 6 nsew
flabel metal1 1430 -4000 1630 -3800 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
