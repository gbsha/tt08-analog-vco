magic
tech sky130A
timestamp 1725567059
<< metal1 >>
rect -1300 3635 -555 3735
rect 2735 3635 2995 3735
rect 6285 3635 7005 3740
rect -1300 -4975 -1200 3635
rect 795 3155 895 3255
rect 1285 3155 1385 3255
rect 4345 3155 4445 3255
rect 4835 3155 4935 3255
rect -1125 2795 -555 2830
rect -1125 -400 -1055 2795
rect 2735 2765 2995 2865
rect 6285 2795 6830 2830
rect 6285 2125 6705 2185
rect 2655 1330 2715 2115
rect 2655 1280 3075 1330
rect -990 625 -455 630
rect -990 585 -550 625
rect -1140 -500 -1040 -400
rect -1125 -4135 -1055 -500
rect -990 -3485 -920 585
rect -555 535 -550 585
rect -460 535 -455 625
rect -555 530 -455 535
rect -850 430 -555 490
rect 3015 465 3075 1280
rect -850 -1670 -780 430
rect 6290 330 6580 390
rect 2635 270 2735 290
rect 2635 265 2900 270
rect 2635 230 2835 265
rect 2735 210 2835 230
rect 2830 135 2835 210
rect 2895 135 2900 265
rect 2830 130 2900 135
rect -705 -500 -555 -400
rect 2735 -500 2995 -400
rect 6285 -500 6450 -400
rect -705 -840 -605 -500
rect -510 -715 -410 -615
rect 2735 -770 2995 -570
rect -705 -940 -555 -840
rect 2735 -940 2995 -840
rect 6285 -940 6450 -840
rect 2830 -1475 2900 -1470
rect 2830 -1605 2835 -1475
rect 2895 -1550 2900 -1475
rect 2895 -1605 2995 -1550
rect 2830 -1610 2995 -1605
rect 6505 -1635 6580 330
rect -850 -1730 -560 -1670
rect 6505 -1725 6510 -1635
rect 6575 -1725 6580 -1635
rect 6505 -1730 6580 -1725
rect 6635 -1770 6705 2125
rect 6145 -1830 6705 -1770
rect 2655 -2620 2715 -1850
rect 2655 -2670 3075 -2620
rect 3015 -3455 3075 -2670
rect -990 -3535 -555 -3485
rect -990 -3540 -705 -3535
rect -1125 -4170 -555 -4135
rect 2735 -4205 2995 -4105
rect 6790 -4135 6830 2795
rect 6285 -4170 6830 -4135
rect 795 -4595 895 -4495
rect 1285 -4595 1385 -4495
rect 4345 -4595 4445 -4495
rect 4835 -4595 4935 -4495
rect 6890 -4975 7005 3635
rect -1300 -5075 -555 -4975
rect 2735 -5075 2995 -4975
rect 6285 -5075 7005 -4975
<< via1 >>
rect -550 535 -460 625
rect 2835 135 2895 265
rect 2835 -1605 2895 -1475
rect 6510 -1725 6575 -1635
<< metal2 >>
rect -555 625 -455 630
rect -555 535 -550 625
rect -460 535 -455 625
rect -555 530 -455 535
rect 2830 265 2900 270
rect 2830 135 2835 265
rect 2895 135 2900 265
rect 2830 130 2900 135
rect 2830 -1475 2900 -1470
rect 2830 -1605 2835 -1475
rect 2895 -1605 2900 -1475
rect 2830 -1610 2900 -1605
rect 6505 -1635 6580 -1630
rect 6505 -1725 6510 -1635
rect 6575 -1725 6580 -1635
rect 6505 -1730 6580 -1725
<< via2 >>
rect -550 535 -460 625
rect 2835 135 2895 265
rect 2835 -1605 2895 -1475
rect 6510 -1725 6575 -1635
<< metal3 >>
rect -555 625 -455 630
rect -555 535 -550 625
rect -460 535 -455 625
rect -555 530 -455 535
rect 2830 265 2900 270
rect 2830 135 2835 265
rect 2895 135 2900 265
rect 2830 130 2900 135
rect 2830 -1475 2900 -1470
rect 2830 -1605 2835 -1475
rect 2895 -1605 2900 -1475
rect 2830 -1610 2900 -1605
rect 6505 -1635 6580 -1630
rect 6505 -1725 6510 -1635
rect 6575 -1725 6580 -1635
rect 6505 -1730 6580 -1725
<< via3 >>
rect -550 535 -460 625
rect 2835 135 2895 265
rect 2835 -1605 2895 -1475
rect 6510 -1725 6575 -1635
<< metal4 >>
rect -555 625 -455 630
rect -555 535 -550 625
rect -460 535 -455 625
rect -555 530 -455 535
rect 2830 265 2900 270
rect 2830 135 2835 265
rect 2895 190 2900 265
rect 2895 135 2995 190
rect 2830 130 2995 135
rect 2735 -1475 2900 -1470
rect 2735 -1530 2835 -1475
rect 2830 -1605 2835 -1530
rect 2895 -1605 2900 -1475
rect 2830 -1610 2900 -1605
rect 6505 -1635 6580 -1630
rect 6505 -1725 6510 -1635
rect 6575 -1725 6580 -1635
rect 6505 -1870 6580 -1725
rect 6185 -1925 6580 -1870
use vco_stage  x1
timestamp 1725560742
transform 1 0 -1400 0 1 980
box 840 -1650 4135 2760
use vco_stage  x2
timestamp 1725560742
transform -1 0 7130 0 1 980
box 840 -1650 4135 2760
use vco_stage  x3
timestamp 1725560742
transform -1 0 7130 0 -1 -2320
box 840 -1650 4135 2760
use vco_stage  x4
timestamp 1725560742
transform 1 0 -1400 0 -1 -2320
box 840 -1650 4135 2760
<< labels >>
flabel metal1 -510 -715 -410 -615 0 FreeSans 128 0 0 0 VSS
port 1 nsew
flabel metal1 -705 -720 -605 -620 0 FreeSans 128 0 0 0 Vc
port 3 nsew
flabel metal1 -1300 3635 -1200 3735 0 FreeSans 128 0 0 0 VDD
port 0 nsew
flabel metal1 -1140 -500 -1040 -400 0 FreeSans 128 0 0 0 Vb
port 2 nsew
flabel metal1 795 3155 895 3255 0 FreeSans 128 0 0 0 Vp0
port 4 nsew
flabel metal1 1285 3155 1385 3255 0 FreeSans 128 0 0 0 Vn0
port 8 nsew
flabel metal1 4835 -4595 4935 -4495 0 FreeSans 128 0 0 0 Vp2
port 6 nsew
flabel metal1 4345 -4595 4445 -4495 0 FreeSans 128 0 0 0 Vn2
port 10 nsew
flabel metal1 795 -4595 895 -4495 0 FreeSans 128 0 0 0 Vp3
port 7 nsew
flabel metal1 1285 -4595 1385 -4495 0 FreeSans 128 0 0 0 Vn3
port 11 nsew
flabel metal1 4345 3155 4445 3255 0 FreeSans 128 0 0 0 Vn1
port 9 nsew
flabel metal1 4835 3155 4935 3255 0 FreeSans 128 0 0 0 Vp1
port 5 nsew
<< end >>
