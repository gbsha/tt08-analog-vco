magic
tech sky130A
magscale 1 2
timestamp 1725533225
<< locali >>
rect 4280 -1550 5680 -1320
rect 4280 -2290 4400 -1550
rect 5560 -2290 5680 -1550
rect 4280 -2430 5680 -2290
<< metal1 >>
rect 1690 5320 1890 5520
rect 4390 4350 4590 4550
rect 5370 4350 5570 4550
rect 1690 3570 1890 3770
rect 4830 2960 4940 3460
rect 5120 3320 5130 3520
rect 5330 3320 5340 3520
rect 4830 2830 5130 2960
rect 1690 2270 1890 2470
rect 4620 2260 4630 2460
rect 4830 2260 4840 2460
rect 5020 2330 5130 2830
rect 8070 2270 8270 2470
rect 1690 -1140 1890 -940
rect 8070 -1140 8270 -940
rect 4440 -2560 4500 -1720
rect 4710 -2150 4780 -1650
rect 4940 -1730 5010 -1720
rect 4940 -2120 5010 -2110
rect 5170 -2150 5240 -1650
rect 4560 -2220 4570 -2150
rect 4840 -2220 4850 -2150
rect 5100 -2220 5110 -2150
rect 5380 -2220 5390 -2150
rect 5450 -2560 5510 -1720
rect 1690 -2770 8270 -2760
rect 1690 -2950 4520 -2770
rect 4700 -2950 5250 -2770
rect 5430 -2950 8270 -2770
rect 1690 -2960 8270 -2950
rect 1690 -3300 1890 -3100
<< via1 >>
rect 5130 3320 5330 3520
rect 4630 2260 4830 2460
rect 4940 -2110 5010 -1730
rect 4570 -2220 4840 -2150
rect 5110 -2220 5380 -2150
rect 4520 -2950 4700 -2770
rect 5250 -2950 5430 -2770
<< metal2 >>
rect 5130 3520 5330 3530
rect 5120 3460 5130 3520
rect 5020 3320 5130 3460
rect 5330 3320 5340 3520
rect 5020 3310 5330 3320
rect 5020 2960 5130 3310
rect 4830 2830 5130 2960
rect 4830 2470 4940 2830
rect 4630 2460 4940 2470
rect 4830 2330 4940 2460
rect 4630 2250 4830 2260
rect 4940 -1730 5010 -1720
rect 4560 -2220 4570 -2150
rect 4840 -2220 4850 -2150
rect 4560 -2760 4660 -2220
rect 4510 -2770 4710 -2760
rect 4510 -2950 4520 -2770
rect 4700 -2950 4710 -2770
rect 4510 -2960 4710 -2950
rect 4940 -3100 5010 -2110
rect 5100 -2220 5110 -2150
rect 5380 -2220 5390 -2150
rect 5290 -2760 5390 -2220
rect 5240 -2770 5440 -2760
rect 5240 -2950 5250 -2770
rect 5430 -2950 5440 -2770
rect 5240 -2960 5440 -2950
rect 4690 -3300 5270 -3100
use sky130_fd_pr__nfet_01v8_XVWV9B  sky130_fd_pr__nfet_01v8_XVWV9B_1
timestamp 1725469944
transform 1 0 4975 0 1 -1920
box -625 -410 625 410
use vco_stage_half  vco_stage_half_0
timestamp 1725531458
transform 1 0 260 0 1 2060
box 1430 -5360 4720 3450
use vco_stage_half  vco_stage_half_1
timestamp 1725531458
transform -1 0 9700 0 1 2060
box 1430 -5360 4720 3450
<< labels >>
flabel metal1 4390 4350 4590 4550 0 FreeSans 1280 0 0 0 Vpbuf
port 8 nsew
flabel metal1 5370 4350 5570 4550 0 FreeSans 1280 0 0 0 Vnbuf
port 9 nsew
flabel metal1 1690 5320 1890 5520 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 1690 -3300 1890 -3100 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 1690 -2960 1890 -2760 0 FreeSans 1280 0 0 0 Vc
port 5 nsew
flabel metal1 1690 -1140 1890 -940 0 FreeSans 1280 0 0 0 Vp
port 2 nsew
flabel metal1 1690 3570 1890 3770 0 FreeSans 1280 0 0 0 Vb
port 4 nsew
flabel metal1 1690 2270 1890 2470 0 FreeSans 1280 0 0 0 Vpout
port 6 nsew
flabel metal1 8070 2270 8270 2470 0 FreeSans 1280 0 0 0 Vnout
port 7 nsew
flabel metal1 8070 -1140 8270 -940 0 FreeSans 1280 0 0 0 Vn
port 3 nsew
<< end >>
