** sch_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_core.sch
.subckt vco_core VDD VSS Vb Vc Vp0 Vp1 Vp2 Vp3 Vn0 Vn1 Vn2 Vn3
*.PININFO VDD:B VSS:B Vb:I Vc:I Vp0:O Vp1:O Vp2:O Vp3:O Vn0:O Vn1:O Vn2:O Vn3:O
x1 VDD VSS Vp Vn Vb Vc net1 net2 Vp0 Vn0 vco_stage
x2 VDD VSS net1 net2 Vb Vc net3 net4 Vp1 Vn1 vco_stage
x3 VDD VSS net3 net4 Vb Vc net5 net6 Vp2 Vn2 vco_stage
x4 VDD VSS net5 net6 Vb Vc Vn Vp Vp3 Vn3 vco_stage
.ends

* expanding   symbol:  vco_stage.sym # of pins=10
** sym_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_stage.sym
** sch_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_stage.sch
.subckt vco_stage VDD VSS Vp Vn Vb Vc Vpout Vnout Vpbuf Vnbuf
*.PININFO VDD:B VSS:B Vp:I Vn:I Vb:I Vc:I Vpout:O Vnout:O Vpbuf:O Vnbuf:O
x1 VDD VSS Vp Vb Vnout Vpout Vds_m5 Vpbuf vco_stage_half
x2 VDD VSS Vn Vb Vpout Vnout Vds_m5 Vnbuf vco_stage_half
XM5 Vds_m5 Vc VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=4 nf=2 m=1
.ends


* expanding   symbol:  vco_stage_half.sym # of pins=8
** sym_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_stage_half.sym
** sch_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_stage_half.sch
.subckt vco_stage_half VDD VSS Vin Vb Vd Vout Vs Vbuf
*.PININFO VDD:B VSS:B Vin:I Vb:I Vd:I Vout:O Vs:O Vbuf:O
XM7 Vout Vd VDD VDD sky130_fd_pr__pfet_01v8 L=2 W=4 nf=2 m=1
XM3 Vout Vb VDD VDD sky130_fd_pr__pfet_01v8 L=2 W=4 nf=2 m=1
XM1 Vout Vin Vs VSS sky130_fd_pr__nfet_01v8 L=2 W=4 nf=2 m=1
x1 VDD VSS Vout Vbuf vco_buffer
XM8 VSS Vout VSS VSS sky130_fd_pr__nfet_01v8 L=11 W=11 nf=1 m=1
.ends


* expanding   symbol:  vco_buffer.sym # of pins=4
** sym_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_buffer.sym
** sch_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_buffer.sch
.subckt vco_buffer VDD VSS Vin Vout
*.PININFO VDD:B VSS:B Vin:I Vout:O
x1 VDD Vin net1 VSS vco_inverter
x2 VDD net1 Vout VSS vco_inverter
.ends


* expanding   symbol:  vco_inverter.sym # of pins=4
** sym_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_inverter.sym
** sch_path: /foss/designs/git/gbsha/tt08-analog-vco/xschem/vco_inverter.sch
.subckt vco_inverter VDD Vin Vout VSS
*.PININFO VDD:B VSS:B Vin:I Vout:O
XM1 Vout Vin VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
